-- File:	WOKBuilder_MSHeaderExtractor.cdl
-- Created:	Tue Mar 19 19:26:26 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1996


class    MSHeaderExtractor from WOKBuilder 
inherits MSExtractor     from WOKBuilder 

	---Purpose: 

uses
    MSActionStatus          from WOKBuilder,
    MSActionType            from WOKBuilder,
    MSAction                from WOKBuilder,
    Param                   from WOKUtils,
    TimeStat                from WOKUtils,
    HAsciiString            from TCollection,
    HSequenceOfHAsciiString from TColStd

is
    
    Create(ashared    : HAsciiString from TCollection;
    	   searchlist : HSequenceOfHAsciiString from TColStd)
    	returns mutable MSHeaderExtractor from WOKBuilder;
    
    Create (
     aname      : HAsciiString            from TCollection;
     ashared    : HAsciiString            from TCollection;
     searchlist : HSequenceOfHAsciiString from TColStd
    ) returns mutable MSHeaderExtractor from WOKBuilder;

    Create(aname : HAsciiString from TCollection; params : Param from WOKUtils)
    	returns mutable MSHeaderExtractor from WOKBuilder;

    Create(params : Param from WOKUtils) 
    	returns mutable MSHeaderExtractor from WOKBuilder;

    GetTypeDepList(me; atype : HAsciiString from TCollection)
    	returns HSequenceOfHAsciiString from TColStd
	is protected;

    GetTypeMDate(me;  atype : HAsciiString from TCollection)
    	returns TimeStat from WOKUtils;
    
    ExtractorID(me)
    	returns MSActionType from WOKBuilder
    	is redefined;

    ExtractionStatus(me:mutable; anaction : MSAction from WOKBuilder)
    	returns MSActionStatus from WOKBuilder
    	is redefined;

end MSHeaderExtractor;
