-- File:	WOKMake_OutputFile.cdl
-- Created:	Thu Apr 25 21:54:16 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1996


class    OutputFile from WOKMake 
inherits StepFile   from WOKMake

	---Purpose: 

uses
    Locator                                  from WOKernel,
    File                                     from WOKernel,
    Entity                                   from WOKBuilder,
    IndexedDataMapOfHAsciiStringOfOutputFile from WOKMake,
    HSequenceOfOutputFile                    from WOKMake,
    FileStatus                               from WOKMake,
    InputFile                                from WOKMake,
    Path                                     from WOKUtils,
    HAsciiString                             from TCollection

is

    Create returns mutable OutputFile  from WOKMake;

    Create(anid      : HAsciiString from TCollection;
    	   afile     : File from WOKernel; 
           abuildent : Entity from WOKBuilder; 
           aoldpath  : Path from WOKUtils)
    	returns mutable OutputFile  from WOKMake;

    Create(aninfile : InputFile from WOKMake)
    	returns mutable OutputFile from WOKMake;
	
    --
    --     READ/WRITE OUTPUT FILES 
    --  

    ReadLine(myclass; astream     : out IStream from Standard;
    	    	      locator     : Locator from WOKernel;
    	    	      infile      : out OutputFile from WOKMake)
    	is private;

    WriteLine(myclass; astream     : out OStream from Standard;
    	    	       infile      : OutputFile from WOKMake)
        is private;

    -- Into/From a map
    ReadFile(myclass;    afile : Path from WOKUtils; 
    	    	      alocator : Locator from WOKernel;
    	    	          amap : out IndexedDataMapOfHAsciiStringOfOutputFile from WOKMake)
    	returns Integer from Standard;
    
    WriteFile(myclass; afile : Path from WOKUtils; amap : IndexedDataMapOfHAsciiStringOfOutputFile from WOKMake)
    	returns Integer from Standard;
	
    -- Into/From a seq
    ReadFile(myclass; afile    : Path from WOKUtils; 
    	    	      alocator : Locator from WOKernel;
    	    	      aseq     : HSequenceOfOutputFile from WOKMake)
    	returns Integer from Standard;
    
    WriteFile(myclass; afile : Path from WOKUtils; aseq : HSequenceOfOutputFile from WOKMake)
    	returns Integer from Standard;

    SetReference(me:mutable);
    SetProduction(me:mutable);
    
    IsProduction(me) returns Boolean from Standard;
    ---C++: inline
     
    SetMember(me:mutable);
    SetExtern(me:mutable);
     
    IsMember(me) 
    ---C++: inline
    	returns Boolean from Standard;

end OutputFile;
