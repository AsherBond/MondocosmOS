-- File:	WOKStep_EngineExtract.cdl
-- Created:	Thu Jun 27 17:22:16 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class EngineExtract from WOKStep 
inherits Extract from WOKStep

	---Purpose: 

uses
    BuildProcess          from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    InputFile             from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection
 
is

    Create(abp   : BuildProcess    from WOKMake; 
    	   aunit : DevUnit         from WOKernel; 
    	   acode : HAsciiString    from TCollection; 
    	   checked, hidden : Boolean  from Standard) 
    	returns mutable EngineExtract from WOKStep;

    HandleInputFile(me:mutable; item : InputFile from WOKMake) 
    	returns Boolean from Standard
    	is redefined protected;

    OutOfDateEntities(me:mutable) 
    	returns HSequenceOfInputFile from WOKMake
    	is redefined protected;
    
end EngineExtract;
