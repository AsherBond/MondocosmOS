-- File:	MS_Engine.cdl
-- Created:	Mon Aug 23 18:19:49 1993
-- Author:	Christophe LEYNADIER
--		<cle@ilebon>
---Copyright:	 Matra Datavision 1993

class Engine 
	---Purpose: 

    from 
    	MS 
    inherits Exec from MS 
    uses 
    	HSequenceOfHAsciiString from TColStd,
	HAsciiString from TCollection

is

    Create(anEngine :HAsciiString) 
    	returns mutable Engine from MS;
    
    Use(me: mutable; aEngine: HAsciiString);
    Uses(me) returns mutable HSequenceOfHAsciiString from TColStd;
          
    Interface(me: mutable; aInterface: HAsciiString);
    Interfaces(me) returns mutable HSequenceOfHAsciiString from TColStd;

fields

    myUses       : HSequenceOfHAsciiString from TColStd;
    myInterfaces : HSequenceOfHAsciiString from TColStd;

end Engine from MS;


