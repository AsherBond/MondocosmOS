-- File:	MSAPI_MemberMet.cdl
-- Created:	Tue Sep 19 22:13:54 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class MemberMet from MSAPI 

	---Purpose: 

uses
    ArgTable     from WOKTools,
    Return       from WOKTools
is

    Info(myclass; argc : Integer from Standard; argv : ArgTable from WOKTools; values : out Return from WOKTools) 
    	returns Integer from Standard;

end MemberMet;
