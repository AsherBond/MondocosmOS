-- File:	WOKBuilder_ImportLibrary.cdl
-- Created:	Wed Oct 23 09:29:38 1996
-- Author:	PLOTNIKOV Eugeny
--		<eugeny@maniax>
---Copyright:	 Matra Datavision 1996

class ImportLibrary from WOKBuilder inherits Library from WOKBuilder

 uses
    
    Path             from WOKUtils, 
    Param            from WOKUtils,
    LibReferenceType from WOKBuilder,
    HAsciiString     from TCollection

 is

    Create (apth  : Path from WOKUtils ) 
     returns mutable ImportLibrary from WOKBuilder;

    Create (
     aname    : HAsciiString     from TCollection; 
     adir     : Path             from WOKUtils; 
     areftype : LibReferenceType from WOKBuilder
    ) returns mutable ImportLibrary from WOKBuilder;

    GetLibFileName (
     me     : mutable;
     params : Param  from  WOKUtils
    ) returns HAsciiString from TCollection is redefined static;
  
    GetLibFileName (
     myclass;
     params : Param        from  WOKUtils;
     aname  : HAsciiString from TCollection
    ) returns HAsciiString from TCollection;

end ImportLibrary;
