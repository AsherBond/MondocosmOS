-- File:	WOKStep_Source.cdl
-- Created:	Thu Jun 27 17:15:36 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class Source from WOKStep 
inherits Step from WOKMake

	---Purpose: Computes Source File List.

uses
    BuildProcess         from WOKMake,
    InputFile            from WOKMake,
    HSequenceOfInputFile from WOKMake,
    DevUnit              from WOKernel,
    File                 from WOKernel,
    HSequenceOfFile      from WOKernel,
    HSequenceOfEntity    from WOKBuilder,
    HAsciiString         from TCollection

is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel; 
    	   acode    : HAsciiString    from TCollection;
    	   checked, hidden : Boolean  from Standard)  
    	returns mutable Source from WOKStep;

    AdmFileType(me)
    	returns HAsciiString from TCollection
        is redefined protected;
    
    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;
    
    HandleInputFile(me:mutable; anitem : InputFile from WOKMake)
    	returns Boolean from Standard
    	is redefined protected;

    GetFILES(me) 
    	returns File from WOKernel
    	is  protected;

    ReadFILES(me:mutable; FILES : InputFile from WOKMake) 
    	is virtual protected;
    
    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake)
    ---Purpose: Executes step    
    --          Computes output files
    	is redefined private;


end Source;
