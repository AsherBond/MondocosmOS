-- File:	WOKStep_SourceExtract.cdl
-- Created:	Thu Jun 27 17:21:38 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class SourceExtract from WOKStep
inherits Extract from WOKStep

	---Purpose: 

uses
    BuildProcess          from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection

is
    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel;
    	   acode    : HAsciiString    from TCollection; 
    	   checked, hidden : Boolean  from Standard) 
    	returns mutable SourceExtract from WOKStep;

    AdmFileType(me)
    	returns HAsciiString from TCollection
        is redefined protected;

    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

    OutOfDateEntities(me:mutable) 
    ---Purpose: Set Build flag to OutOfDate entities 
    --          Clears Build flag to Uptodate Entities
    --          This base implementation does nothing
    	returns HSequenceOfInputFile from WOKMake
    	is redefined protected;

    
    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake) 
    	is redefined private;

end SourceExtract;
