-- File:	WOKTools_CStringHasher.cdl
-- Created:	Fri Jul 19 16:28:16 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class CStringHasher from WOKTools
uses
    CString from Standard
is

   HashCode(myclass; Key : CString from Standard) returns Integer;
	    ---Level: Public
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	-- range 0..Upper.
	-- Default ::HashCode(K,Upper)
	    
   IsEqual(myclass; K1, K2 : CString from Standard) returns Boolean;
	---Level: Public
	---Purpose: Returns True  when the two  keys are the same. Two
	-- same  keys  must   have  the  same  hashcode,  the
	-- contrary is not necessary.
	-- Default K1 == K2
end;
