-- File:	WOKUnix_Buffer.cdl
-- Created:	Thu May  4 16:33:47 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995

private deferred class Buffer from WOKUnix
inherits TShared from MMgt
uses 
    BufferIs from WOKUnix,
    FDescr   from WOKUnix,
    FDSet    from WOKUnix,
    Timeval  from WOKUnix,
    HSequenceOfHAsciiString from TColStd
    
raises
    BufferOverflow from WOKUnix,
    ProcessTimeOut from WOKUnix
is
    Initialize(afd : FDescr   from WOKUnix; astd : BufferIs from WOKUnix);

    Clear(me : mutable);
    
    GetFDescr(me) returns FDescr from WOKUnix;
    SetFDescr(me:mutable; afd : FDescr from WOKUnix);

    BufferIs(me) returns BufferIs from WOKUnix;  
    AssociatedChannel(me) returns FDescr from WOKUnix;
    
    Select(me; afd : out Integer; atimeout : in out Timeval from WOKUnix; aset : in out FDSet from WOKUnix) is deferred;
    Acquit(me:mutable;  astatus : Integer from Standard; aset : FDSet from WOKUnix) raises ProcessTimeOut from WOKUnix is deferred;
    
    Echo(me : mutable)   returns HSequenceOfHAsciiString from TColStd is virtual;
    Errors(me : mutable) returns HSequenceOfHAsciiString from TColStd is virtual;
 
    Write(me : mutable ; afd : in out FDescr from WOKUnix) ;
    
    Close(me:mutable) is virtual;
    
fields
    myfd  : FDescr from WOKUnix;
    mystd : BufferIs from WOKUnix;
end;
