-- File:	WOKTCL.cdl
-- Created:	Fri Aug 11 11:33:51 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


package WOKTCL 

	---Purpose: 

uses 
    
    WOKTclTools,
    WOKTools,
    WOKAPI

is

    class Interpretor;

    ---class LocatorTable
    ---	instantiates HandleTable from WOKTclTools ( Locator from WOKAPI );

end WOKTCL;
