-- File:	WOKDeliv_DeliverySTUBClient.cdl
-- Created:	Mon Aug 19 11:37:28 1996
-- Author:	Arnaud BOUZY
--		<adn@legox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class DeliverySTUBClient from WOKDeliv inherits DeliveryMetaStep from WOKDeliv

	---Purpose: Process interfaces for delivery units (client stub) 

uses DevUnit from WOKernel,
     File from WOKernel,
     BuildProcess from WOKMake,
     InputFile from WOKMake,
     HSequenceOfInputFile from WOKMake,
     HAsciiString from TCollection

is

    Create(abp      : BuildProcess from WOKMake;
    	   aunit    : DevUnit from WOKernel; 
    	   acode    : HAsciiString from TCollection; 
    	   checked, hidden : Boolean  from Standard)
    returns mutable DeliverySTUBClient from WOKDeliv;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake)
    is private;
    
    HandleInputFile(me:mutable; anitem : InputFile from WOKMake)
    returns Boolean from Standard
    is protected;
    
    AdmFileType(me)
    	returns HAsciiString from TCollection;


end DeliverySTUBClient;
