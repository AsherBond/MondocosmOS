-- File:	WOKernel_Workbench.cdl
-- Created:	Fri Jun 23 17:49:24 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class Workbench from WOKernel 
inherits UnitNesting from WOKernel

	---Purpose: a workbench is the developing Environment of a developper

uses
    HAsciiString                from TCollection,
    Workshop                    from WOKernel,
    FileType                    from WOKernel,
    File                        from WOKernel,
    Locator                     from WOKernel,
    HSequenceOfParamItem        from WOKUtils,
    HSequenceOfHAsciiString     from TColStd

raises
    ProgramError from Standard
is

    Create(aname : HAsciiString from TCollection; anesting : Workshop from WOKernel; afather : Workbench from WOKernel)   
    ---Purpose: Instantiates a workbench    
    	returns mutable Workbench from  WOKernel; 
    
    GetParameters(me:mutable)
    is redefined protected;

    EntityCode(me) 
    	returns HAsciiString from TCollection
	is redefined;

    GetUnitList(me:mutable)
    	returns HSequenceOfHAsciiString from TColStd
	is redefined private;

    GetUnitListFile(me)
    	returns File from WOKernel
	is redefined private;

    Open(me: mutable)
    ---Purpose: Opens an existing Workbench    
    	raises ProgramError from Standard is redefined; 
	
    Close(me: mutable) is redefined;
    ---Purpose: Closes an Opened Workbench
     
    Father(me) returns mutable HAsciiString from TCollection;
    ---Purpose: Gives the Father Workbench of me    
    
    SetFather(me:mutable; afather : Workbench from WOKernel);
    ---Purpose: Set the father of Wb    
    
    Ancestors(me) returns HSequenceOfHAsciiString from TColStd;
    ---Purpose: Gives the ancestors of me

    Visibility(me) returns HSequenceOfHAsciiString from TColStd;
    ---Purpose: Gives The nestings in visibility of workbench    

fields
    myfather     : HAsciiString from TCollection;
end Workbench;
