-- File:	WOKTools_AsciiStringHasher.cdl
-- Created:	Tue May 30 10:03:37 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class AsciiStringHasher from WOKTools
uses
    AsciiString from TCollection
is

   HashCode(myclass; Key : AsciiString from TCollection) returns Integer;
	    ---Level: Public
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	-- range 0..Upper.
	-- Default ::HashCode(K,Upper)
	    
   IsEqual(myclass; K1, K2 : AsciiString from TCollection) returns Boolean;
	---Level: Public
	---Purpose: Returns True  when the two  keys are the same. Two
	-- same  keys  must   have  the  same  hashcode,  the
	-- contrary is not necessary.
	-- Default K1 == K2
end;
