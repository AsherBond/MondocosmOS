-- File:	WOKDFLT_DFLTExtract.cdl
-- Created:	Fri Jun  7 11:21:39 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class DFLTExtract from WOKDFLT 
inherits Extract from WOKStep

	---Purpose: 

uses
    BuildProcess          from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection

is

    Create(abp   : BuildProcess from WOKMake;
    	   aunit : DevUnit from WOKernel; 
    	   acode : HAsciiString from TCollection;
    	   checked, hidden : Boolean  from Standard) 
    	returns mutable DFLTExtract from WOKDFLT;

    OutOfDateEntities(me:mutable) 
    	returns HSequenceOfInputFile from WOKMake
    	is redefined protected;

end DFLTExtract;
