-- File:	WOKStep_ExtractExecList.cdl
-- Created:	Wed Aug 28 18:22:45 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class ExtractExecList from WOKStep 
inherits     MetaStep from WOKMake

	---Purpose: 

uses
    BuildProcess            from WOKMake,
    HSequenceOfInputFile    from WOKMake,
    InputFile               from WOKMake,
    DevUnit                 from WOKernel,
    HSequenceOfHAsciiString from TColStd,
    HAsciiString            from TCollection

is
    Create( abp      : BuildProcess    from WOKMake; 
    	    aunit    : DevUnit         from WOKernel; 
    	    acode    : HAsciiString    from TCollection; 
    	    checked, hidden : Boolean  from Standard)
    	returns mutable ExtractExecList from WOKStep;
	       
    HandleInputFile(me:mutable; anitem : InputFile from WOKMake)
    	returns Boolean from Standard
    	is redefined protected;

    AdmFileType(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake) 
    ---Purpose: Executes underlying steps
    --          Computes output files
    	is redefined private;

end ExtractExecList;
