-- File:	WOKBuilder_DLLFile.cdl
-- Created:	Mon Oct 21 14:10:20 1996
-- Author:	PLOTNIKOV Eugeny
--		<eugeny@maniax>
---Copyright:	 Matra Datavision 1996

class DLLFile from WOKBuilder inherits Entity  from WOKBuilder 

 uses
    
    Path from WOKUtils

 is

    Create ( apath : Path from WOKUtils ) returns mutable DLLFile from WOKBuilder;

end DLLFile;
