
-- -- File:	WOKernel_UnitNesting.cdl
-- Created:	Fri Jun 23 18:31:37 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


deferred class UnitNesting from WOKernel 
inherits Entity from WOKernel

	---Purpose: 

uses
    Entity                  from WOKernel,
    DevUnit                 from WOKernel,
    HSequenceOfDBMSID       from WOKernel,
    HSequenceOfStationID    from WOKernel,
    UnitTypeBase            from WOKernel,
    FileType                from WOKernel,
    FileTypeBase            from WOKernel,
    File                    from WOKernel,
    Path                    from WOKUtils,
    HSequenceOfParamItem    from WOKUtils,
    HAsciiString            from TCollection,
    HSequenceOfHAsciiString from TColStd

raises
    ProgramError from Standard
is
    Initialize(aname : HAsciiString from TCollection; anesting : Entity from WOKernel);

    GetUnitList(me:mutable)
    	returns HSequenceOfHAsciiString from TColStd
	is deferred private;

    GetUnitListFile(me)
    	returns File from WOKernel
	is deferred private;

    Open(me: mutable)  
    	raises ProgramError from Standard;

    Close(me: mutable);
   
    Units(me) 
    	returns HSequenceOfHAsciiString from TColStd is static;

    DumpUnitList(me) is static private;

    GetDevUnit(me; akey : Character from Standard; aname : HAsciiString from TCollection)
    	returns DevUnit from WOKernel;
	
    GetDevUnit(me; atype, aname : HAsciiString from TCollection)
    	returns DevUnit from WOKernel;

    KnownTypes(me) 
    ---C++: return const &
       	returns UnitTypeBase from WOKernel;

    AddUnit(me:mutable; aunit : DevUnit from WOKernel) 
    	raises ProgramError from Standard is static;

    RemoveUnit(me:mutable; aunit : DevUnit from WOKernel) 
    	raises ProgramError from Standard is static;

fields
    mytypebase : UnitTypeBase                  from WOKernel;
    myunits    : HSequenceOfHAsciiString       from TColStd;
end UnitNesting;
