-- File:	WOKStep_TransitiveLinkList.cdl
-- Created:	Tue Dec  2 18:16:48 1997
-- Author:	Jean GAUTIER
--		<jga@hourax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class TransitiveLinkList from WOKStep 
inherits ComputeLinkList from WOKStep

	---Purpose: 

uses
    BuildProcess from WOKMake,
    DevUnit from WOKernel,
    HSequenceOfHAsciiString from TColStd,
    HAsciiString from TCollection

is

    Create( abp      : BuildProcess     from WOKMake; 
    	    aunit    : DevUnit          from WOKernel; 
    	    acode    : HAsciiString     from TCollection; 
    	    checked, hidden : Boolean   from Standard)
    	returns mutable TransitiveLinkList from WOKStep;
 
 
   ComputeDependency(me; code : HAsciiString from TCollection; adirectlist : HSequenceOfHAsciiString from TColStd)
    	returns HSequenceOfHAsciiString from TColStd is redefined protected;

end TransitiveLinkList;
