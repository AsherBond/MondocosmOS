-- File:	WOKBuilder_ObjectFile.cdl
-- Created:	Tue Aug 29 11:26:32 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class ObjectFile from WOKBuilder 
inherits Entity  from WOKBuilder 
	---Purpose: 

uses
    Path from WOKUtils
is

    Create(apath : Path from WOKUtils) returns mutable ObjectFile from WOKBuilder;


end ObjectFile;
