-- File:	WOKOrbix_IDLFill.cdl
-- Created:	Mon Aug 25 11:35:36 1997
-- Author:	Jean GAUTIER
--		<jga@hourax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class IDLFill from WOKOrbix 
inherits Step from WOKMake

	---Purpose: 

uses
    BuildProcess from WOKMake,
    InputFile    from WOKMake,
    HSequenceOfInputFile from WOKMake,
    DevUnit      from WOKernel,
    File         from WOKernel,
    Entity       from WOKBuilder,
    HAsciiString from TCollection

is
    
    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel; 
    	   acode    : HAsciiString    from TCollection; 
    	   checked, hidden : Boolean  from Standard)
    	returns mutable IDLFill from WOKOrbix;

    
    AdmFileType(me)
    	returns HAsciiString from TCollection
        is redefined protected;

    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

    HandleInputFile(me:mutable; item : InputFile from WOKMake) 
    	returns Boolean from Standard
    	is redefined protected;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake) 
    	is redefined private;

end IDLFill;
