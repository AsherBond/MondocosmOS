-- File:	WOKBuilder_CDLFile.cdl
-- Created:	Thu Aug 10 20:49:17 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class CDLFile from WOKBuilder 
inherits Specification from WOKBuilder

	---Purpose: 

uses
    Path from WOKUtils

is

    Create(apath : Path from WOKUtils) returns mutable CDLFile from WOKBuilder;
    
end CDLFile;
