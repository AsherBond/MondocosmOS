-- File:	WOKStep_Library.cdl
-- Created:	Thu Jun 27 17:27:50 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

deferred class Library from WOKStep
inherits Step     from WOKMake

    ---Purpose: 

uses
    BuildProcess          from WOKMake,
    InputFile             from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection
is
    Initialize(abp      : BuildProcess    from WOKMake; 
    	       aunit    : DevUnit         from WOKernel;
    	       acode    : HAsciiString    from TCollection; 
    	       checked, hidden : Boolean  from Standard);

    AdmFileType(me)
    	returns HAsciiString from TCollection
        is redefined protected;

    HandleInputFile(me:mutable; item : InputFile from WOKMake) 
    	returns Boolean from Standard
    	is redefined protected;
	
    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;
   
    CompleteExecList(me:mutable; anexeclist : HSequenceOfInputFile from WOKMake)
    	is redefined protected;

end Library;
