-- File:	WOKStep_DLLink.cdl
-- Created:	Wed Oct 23 10:15:56 1996
-- Author:	PLOTNIKOV Eugeny
--		<eugeny@maniax>
---Copyright:	 Matra Datavision 1996

class DLLink from WOKStep inherits WNTLink from WOKStep

 uses
    BuildProcess            from WOKMake,
    DevUnit                 from WOKernel,
    HAsciiString            from TCollection,
    HSequenceOfLibrary      from WOKBuilder,
    HSequenceOfHAsciiString from TColStd,
    HSequenceOfInputFile    from WOKMake,
    WNTCollector            from WOKBuilder
 
 is
 
    Create (
     aBP     : BuildProcess from WOKMake; 
     aUnit   : DevUnit      from WOKernel;
     aCode   : HAsciiString from TCollection;
     checked : Boolean      from Standard;
     hidden  : Boolean      from Standard
    ) returns mutable DLLink from WOKStep;
    	---Purpose: creates a class instance   

    ComputeLibraryList (
     me      : mutable;
     anInput : HSequenceOfInputFile from WOKMake
    )
     returns mutable HSequenceOfLibrary from WOKBuilder
     is redefined static protected;
     	---Purpose: computes library list to build a target

    ComputeTool ( me : mutable )
     returns mutable WNTCollector from WOKBuilder
     is redefined static protected;
    	---Purpose: computes build tool

end DLLink;
