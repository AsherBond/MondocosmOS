-- File:	WOKTools_BasicMapIterator.cdl
-- Created:	Mon May 29 17:41:11 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995

private deferred class BasicMapIterator from WOKTools 

	---Purpose: This  class  provides    basic   services  for the
	-- iterators  on Maps. The  iterators  are  inherited
	-- from this one.
	-- 
	-- The  iterator   contains  an   array   of pointers
	-- (buckets). Each bucket is a  pointer  on a node. A
	-- node contains a pointer on the next node.
	-- 
	-- This class  provides also basic  services for  the
	-- implementation of Maps.

uses
    BasicMap from WOKTools

is
    Initialize;
	---Purpose: Creates an empty iterator.

    Initialize(M : BasicMap from WOKTools);
	---Purpose: Initialize on the first node in the buckets.
	
    Initialize(me : in out; M : BasicMap from WOKTools)
	---Purpose: Initialize on the first node in the buckets.
    is static protected;
    
    Reset(me : in out)
	---Purpose: Resets the iterator to the first node.
    is static;
    
    More(me) returns Boolean
	---Purpose: Returns True if there is a current  element in the
	--          iterator.
	---C++: inline
    is static;
    
    Next(me : in out)
	---Purpose: Sets the  iterator   to the  next   node.  If  the
	-- iterator is empty it will not change.
    is static;

fields
    	myNbBuckets : Integer;
        myBuckets   : Address from Standard;
        myBucket    : Integer;
        myNode      : Address from Standard is protected;

end BasicMapIterator;
