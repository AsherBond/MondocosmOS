-- File:	WOKernel_Factory.cdl
-- Created:	Fri Jun 23 16:55:29 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class Factory from WOKernel 
inherits Entity from WOKernel


	---Purpose: WOK Factory : corresponds to a developpers Team

uses
    HSequenceOfHAsciiString from TColStd,
    HAsciiString            from TCollection,
    Workshop                from WOKernel,
    Warehouse               from WOKernel,
    Session                 from WOKernel,
    Path                    from WOKUtils,
    HSequenceOfParamItem    from WOKUtils
raises
    ProgramError from Standard
is
    Create(aname : HAsciiString from TCollection; anesting : Session from WOKernel) 
    ---Purpose: instantiates a factory    
    	returns mutable Factory from WOKernel; 
    
    EntityCode(me) 
    	returns HAsciiString from TCollection
	is redefined;

    ReadWSLIST(me:mutable);
    WriteWSList(me:mutable);
    
    Open(me: mutable)
    raises ProgramError from Standard is redefined;
    ---Purpose: opens a factory 
    --          loads Workshop list
    --          load Warehouse parameters
    
    Close(me: mutable) is redefined;
    ---Purpose: closes Factory    

    Workshops(me) 
    ---Purpose: gives the sequence of workshop in factory
    	returns HSequenceOfHAsciiString from TColStd;

    DumpWorkshopList(me);
    ---Purpose: updates files WSLIST with myworkshops    

    AddWorkshop(me:mutable; aworkshop : Workshop from WOKernel)
    ---Purpose: Adds workshop to factory
    --          Updates WSLIST    
    	raises ProgramError from Standard;
   
    RemoveWorkshop(me:mutable; aworkshop : Workshop from WOKernel)
    ---Purpose: removes workshop    
    	raises ProgramError from Standard;
    
    SetWarehouse(me:mutable; awarehouse : Warehouse from WOKernel);
    Warehouse(me) 
    ---Purpose: gives the warehouse of factory    
    	returns HAsciiString from TCollection;
	
    SetSourceStorage(me:mutable; astorage : Path from WOKUtils);
    SourceStorage(me)
    ---Purpose: gives the SCCS repository of factory    
    	returns Path      from WOKUtils;
    
fields
    myworkshops : HSequenceOfHAsciiString from TColStd;
    mywarehouse : HAsciiString            from TCollection;
    mysccsbase  : Path                    from WOKUtils;
end Factory;
