-- File:	WOKStep_ResourceSource.cdl
-- Created:	Thu Sep 26 16:03:25 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


class ResourceSource from WOKStep 
inherits Source from WOKStep 

	---Purpose: 

uses
    BuildProcess from WOKMake,
    DevUnit      from WOKernel,
    InputFile    from WOKMake,
    HAsciiString from TCollection

is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel; 
    	   acode    : HAsciiString    from TCollection;
    	   checked, hidden : Boolean  from Standard)  
    	returns mutable ResourceSource from WOKStep;

    ReadFILES(me:mutable; FILES : InputFile from WOKMake) 
    	is redefined protected;

end ResourceSource;
