-- File:	WOKStep_CDLUnitSource.cdl
-- Created:	Thu Jun 27 17:16:21 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class CDLUnitSource from WOKStep 
inherits Source from WOKStep

	---Purpose: Computes CDLUnitSource File List.

uses
    BuildProcess         from WOKMake,
    HSequenceOfInputFile from WOKMake,
    InputFile            from WOKMake,
    DevUnit              from WOKernel,
    File                 from WOKernel,
    HSequenceOfFile      from WOKernel,
    HSequenceOfEntity    from WOKBuilder,
    HAsciiString         from TCollection

is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel; 
    	   acode    : HAsciiString    from TCollection;  
    	   checked, hidden : Boolean  from Standard)  
    	returns mutable CDLUnitSource from WOKStep;

    GetUnitDescr(me) 
    	returns File from WOKernel
	is protected;

    ReadUnitDescr(me:mutable; unitcdl : InputFile from WOKMake) is virtual protected;
    ---Purpose: Read Unit.cdl file to obtain CDL files list    

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake)
    ---Purpose: Executes step    
    --          Computes output files
    	is redefined private;

end CDLUnitSource;
