-- File:	WOKBuilder_MFile.cdl
-- Created:	Tue Aug 29 11:13:48 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


class MFile from WOKBuilder 
inherits Entity from WOKBuilder

	---Purpose: 

uses
    Path from WOKUtils
is

    Create(apath : Path from WOKUtils) returns mutable MFile from WOKBuilder;


end MFile;
