-- File:	WOKStep_ComputeLinkList.cdl
-- Created:	Tue Sep  3 20:42:48 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996


deferred class ComputeLinkList from WOKStep 
inherits LinkList from WOKStep

	---Purpose: 


uses
    BuildProcess            from WOKMake,
    HSequenceOfInputFile    from WOKMake,
    InputFile               from WOKMake,
    DevUnit                 from WOKernel,
    MapOfHAsciiString       from WOKTools,
    HSequenceOfHAsciiString from TColStd,
    HAsciiString            from TCollection

is

    Initialize( abp      : BuildProcess     from WOKMake; 
    	        aunit    : DevUnit          from WOKernel; 
    	        acode    : HAsciiString     from TCollection; 
    	        checked, hidden : Boolean   from Standard)
    	returns mutable ComputeLinkList from WOKStep;
	       
    HandleInputFile(me:mutable; anitem : InputFile from WOKMake)
    	returns Boolean from Standard
    	is redefined protected;

    AdmFileType(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

    OutputDirTypeName(me)
    	returns HAsciiString from TCollection
    	is redefined protected;

     Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake) 
    	is redefined private;


end ComputeLinkList;
