-- File:	WOKBuilder_Entity.cdl
-- Created:	Thu Aug 10 20:38:52 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


deferred class Entity from WOKBuilder 
inherits TShared from MMgt
	---Purpose: 

uses
    Path              from WOKUtils,
    HSequenceOfEntity from WOKBuilder

raises
    ProgramError from Standard
is
    Initialize(apath : Path from WOKUtils);

    Path(me) 
    ---C++: inline
    ---C++: return const &
       	returns Path from WOKUtils;
    SetPath(me:mutable; apath : Path from WOKUtils);

fields
    mypath       : Path              from WOKUtils;
end Entity;
