-- File:	WOKDeliv_DeliveryOBJSSchema.cdl
-- Created:	Tue Apr 29 10:25:21 1997
-- Author:	Arnaud BOUZY
--		<adn@legox.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class DeliveryOBJSSchema from WOKDeliv inherits DeliveryStep from WOKDeliv

	---Purpose: Process schema for Object Store 

uses DevUnit from WOKernel,
     File from WOKernel,
     BuildProcess from WOKMake,
     InputFile from WOKMake,
     HSequenceOfInputFile from WOKMake,
     HAsciiString from TCollection

is

    Create(aprocess : BuildProcess   from WOKMake;
    	   aunit    : DevUnit from WOKernel; 
    	   acode    : HAsciiString from TCollection; 
    	   checked, hidden : Boolean  from Standard)
    returns mutable DeliveryOBJSSchema from WOKDeliv;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake)
    is private;
    
    HandleInputFile(me:mutable; anitem : InputFile from WOKMake)
    returns Boolean from Standard
    is protected;
    
    AdmFileType(me)
    	returns HAsciiString from TCollection;


end DeliveryOBJSSchema;
