-- File:	WOKStep_DynamicLibrary.cdl
-- Created:	Thu Jun 27 17:30:39 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class DynamicLibrary from WOKStep 
inherits Library from WOKStep

	---Purpose: 

uses
    BuildProcess          from WOKMake,
    InputFile             from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection
is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel;
    	   acode    : HAsciiString    from TCollection; 
    	   checked, hidden : Boolean  from Standard) 
    	returns mutable DynamicLibrary from WOKStep;

    HandleInputFile(me:mutable; item : InputFile from WOKMake) 
    	returns Boolean from Standard
    	is redefined protected;

    ComputeDatabaseDirectories(me)
    	returns HSequenceOfPath from WOKUtils is protected;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake) 
    	is redefined private;

end DynamicLibrary;
