-- File:	WOKAPI_Parcel.cdl
-- Created:	Wed Apr  3 16:40:52 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1996


class Parcel from WOKAPI 
inherits Entity from WOKAPI

	---Purpose: 

uses
    Parcel                  from WOKernel,
    Unit                    from WOKAPI,
    Session                 from WOKAPI,
    Entity                  from WOKAPI,
    SequenceOfUnit          from WOKAPI,
    SequenceOfEntity        from WOKAPI,
    HSequenceOfDefine       from WOKTools,
    HSequenceOfParamItem    from WOKUtils,
    HAsciiString            from TCollection
    
is

    Create returns Parcel from WOKAPI;

    Create(aent : Entity from WOKAPI)
    	returns Parcel from WOKAPI;

    Create(asession : Session from WOKAPI;
    	   aname    : HAsciiString from TCollection;
    	   verbose,getit  : Boolean from Standard = Standard_True)
	returns Parcel from WOKAPI;

    BuildParameters(me; asession : Session from WOKAPI;
    	    	    	apath    : HAsciiString from TCollection;
			defines  : HSequenceOfDefine from WOKTools;
			usedefaults : Boolean from Standard)
    	returns HSequenceOfParamItem from WOKUtils;
    
    Declare(me: in out; asession : Session from WOKAPI;
    	    	    	aname    : HAsciiString from TCollection;
    	    	    	anesting : Entity from WOKAPI;
			defines  : HSequenceOfDefine from WOKTools;
			usedefaults : Boolean from Standard)
    returns Boolean;
    
    Delivery(me; unit : out Unit from WOKAPI);

    NestedEntities(me; aseq : out SequenceOfEntity from WOKAPI)
    	returns Boolean from Standard
    	is redefined;

    Units(me; unitseq : out SequenceOfUnit from WOKAPI);

    IsValid(me) 
    	returns Boolean from Standard
	is redefined;

end Parcel;
