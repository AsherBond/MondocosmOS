-- File:	WOKTools_HAsciiStringHasher.cdl
-- Created:	Wed Jun 28 11:12:13 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995

class HAsciiStringHasher from WOKTools
uses
    HAsciiString from TCollection
is

   HashCode(myclass; Key : HAsciiString from TCollection) returns Integer;
	    ---Level: Public
	---Purpose: Returns a HasCode value  for  the  Key <K>  in the
	-- range 0..Upper.
	-- Default ::HashCode(K,Upper)
	    
   IsEqual(myclass; K1, K2 : HAsciiString from TCollection) returns Boolean;
	---Level: Public
	---Purpose: Returns True  when the two  keys are the same. Two
	-- same  keys  must   have  the  same  hashcode,  the
	-- contrary is not necessary.
	-- Default K1 == K2
end;
