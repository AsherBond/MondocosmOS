-- File:	WOKStep_WNTLibrary.cdl
-- Created:	Fri Oct 25 16:14:54 1996
-- Author:	PLOTNIKOV Eugeny
--		<eugeny@maniax>
---Copyright:	 Matra Datavision 1996

deferred class WNTLibrary from WOKStep inherits WNTCollect from WOKStep

 uses
    BuildProcess         from WOKMake,
    DevUnit              from WOKernel,
    HAsciiString         from TCollection,
    HSequenceOfInputFile from WOKMake,
    InputFile            from WOKMake
    
 is

    Initialize (
     abp     : BuildProcess from WOKMake; 
     aUnit   : DevUnit      from WOKernel;
     aCode   : HAsciiString from TCollection;
     checked : Boolean      from Standard;
     hidden  : Boolean      from Standard
    );
    	---Purpose: provides initialization   
 
    Execute (
     me         : mutable;
     anExecList : HSequenceOfInputFile from WOKMake
    ) is redefined static;
    	---Purpose: executes a tool

    HandleInputFile (
     me     : mutable;
     anItem : InputFile from WOKMake
    ) returns Boolean from Standard is redefined static;
    	---Purpose: adds a file in list if the file is input for step

end WNTLibrary;
