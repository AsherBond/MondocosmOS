-- File:	WOKStep_ClientExtract.cdl
-- Created:	Thu Jun 27 17:20:15 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class ClientExtract from WOKStep 
inherits Extract from WOKStep

	---Purpose: 

uses
    BuildProcess          from WOKMake,
    InputFile             from WOKMake,
    HSequenceOfInputFile  from WOKMake,
    DevUnit               from WOKernel,
    HSequenceOfFile       from WOKernel,
    File                  from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HSequenceOfPath       from WOKUtils,
    HAsciiString          from TCollection
 
is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit         from WOKernel; 
    	   acode    : HAsciiString    from TCollection;
    	   checked, hidden : Boolean  from Standard) 
    	returns mutable ClientExtract from WOKStep;

    HandleInputFile(me:mutable; infile : InputFile from WOKMake)
    	returns Boolean from Standard;

    Init(me:mutable)
    	is redefined protected;

    GetInputFlow(me:mutable)
    	is redefined protected;

    OutOfDateEntities(me:mutable) 
    	returns HSequenceOfInputFile from WOKMake
    	is redefined protected;

    Execute(me:mutable; execlist : HSequenceOfInputFile from WOKMake)
    	is redefined ;

end ClientExtract;
