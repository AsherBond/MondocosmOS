-- File:	WOKStep_ExecutableSource.cdl
-- Created:	Thu Jun 27 17:17:00 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1996

class ExecutableSource from WOKStep
inherits CDLUnitSource from WOKStep

	---Purpose: Computes CDLUnitSource File List.

uses
    BuildProcess          from WOKMake,
    InputFile             from WOKMake,
    DevUnit               from WOKernel,
    File                  from WOKernel,
    HSequenceOfFile       from WOKernel,
    HSequenceOfEntity     from WOKBuilder,
    HAsciiString          from TCollection

is

    Create(abp      : BuildProcess    from WOKMake; 
    	   aunit    : DevUnit from WOKernel; 
    	   acode    : HAsciiString from TCollection;  
    	   checked, hidden : Boolean from Standard)  
    	returns mutable ExecutableSource from WOKStep;

    ReadUnitDescr(me:mutable; unitcdl : InputFile from WOKMake) is redefined protected;
    ---Purpose: Read Unit.cdl file to obtain CDL files list    

end ExecutableSource;


