-- File:	WOKBuilder_MSClientExtractor.cdl
-- Created:	Tue Mar 19 19:32:13 1996
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1996


class MSClientExtractor    from WOKBuilder 
inherits MSHeaderExtractor from WOKBuilder 

	---Purpose: 

uses
    MSActionType            from WOKBuilder,
    MSActionStatus          from WOKBuilder,
    MSAction                from WOKBuilder,
    Param                   from WOKUtils,
    HSequenceOfMemberMet    from MS,
    HSequenceOfExternMet    from MS,
    MapOfHAsciiString       from WOKTools,
    HAsciiString            from TCollection,
    HSequenceOfHAsciiString from TColStd

is

    Create(ashared    : HAsciiString from TCollection;
    	   searchlist : HSequenceOfHAsciiString from TColStd)
    	returns mutable MSClientExtractor from WOKBuilder;
    
    Create(params : Param from WOKUtils) 
    	returns mutable MSClientExtractor from WOKBuilder;

    Init(me:mutable; aname : HAsciiString from TCollection);
    
    MemberMethods(me)
    	returns HSequenceOfMemberMet from MS;
	
    ExternMethods(me)
    	returns HSequenceOfExternMet from MS;
	
    CompleteTypes(me)
    ---C++: return const &
    	returns MapOfHAsciiString    from WOKTools;
    
    IncompleteTypes(me)
    ---C++: return const &
    	returns MapOfHAsciiString    from WOKTools;
    
    SemiCompleteTypes(me)
    ---C++: return const &
    	returns MapOfHAsciiString    from WOKTools;
    
    ExtractorID(me)
    	returns MSActionType from WOKBuilder
    	is redefined;

    ExtractionStatus(me:mutable; anaction : MSAction from WOKBuilder)
    	returns MSActionStatus from WOKBuilder
    	is redefined;

fields

    mycompl  : MapOfHAsciiString    from WOKTools;
    myicompl : MapOfHAsciiString    from WOKTools;
    myscompl : MapOfHAsciiString    from WOKTools;
    mymmeth  : HSequenceOfMemberMet from MS;
    myxmeth  : HSequenceOfExternMet from MS;
    
end MSClientExtractor;
