-- File:	WOKOBJS_LibSchema.cdl
-- Created:	Mon Feb 24 15:04:40 1997
-- Author:	Jean GAUTIER
--		<jga@hourax.paris1.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997


class    LibSchema from WOKOBJS 
inherits Entity    from WOKBuilder

	---Purpose: 

uses
    Path             from WOKUtils, 
    Param            from WOKUtils,
    HAsciiString     from TCollection

is
    
    Create(apth  : Path from WOKUtils) 
    	returns mutable LibSchema from WOKOBJS;

    GetLibFileName(myclass; params : Param  from  WOKUtils; aname : HAsciiString from TCollection) 
    	returns HAsciiString from TCollection;
  

end LibSchema;
